module ctrl_microondas
(
  // Declaração das portas
  //------------
  // COMPLETAR
  //------------
);
	//-----------
	// COMPLETAR
	//-----------
endmodule